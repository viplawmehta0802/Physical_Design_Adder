(*blackbox*)
module four_bit_adder (in1, in2, c_in, out, c_out);
input [3:0] in1, in2;
input c_in;
output [3:0] out;
output c_out;
wire [4:0] sum;

endmodule
